----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    10:15:19 11/25/2021 
-- Design Name: 
-- Module Name:    DeclaracionCaseWhen - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity DeclaracionCaseWhen is port(
A: in std_logic_vector(3 downto 0);
d: out std_logic_vector(6 downto 0));
end DeclaracionCaseWhen;

architecture Behavioral of DeclaracionCaseWhen is
begin
process (A) begin
case A is 
when "0000" = > d < = "0000001"
when "0001" = > d < = "1001111"
when "0010" = > d < = "0010010"
when "0011" = > d < = "0000110"
when "0100" = > d < = "1001100"
when "0101" = > d < = "0100100"
when "0110" = > d < = "0100000"
when "0111" = > d < = "0001110"
when "1000" = > d < = "0000000"
when "1001" = > d < = "0000100"
when others = > d < = "1111111"
end case;
end process;
end Behavioral;

