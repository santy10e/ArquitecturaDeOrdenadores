----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    18:46:55 11/23/2021 
-- Design Name: 
-- Module Name:    WithSelect - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity WithSelect is port(
	a: in std_logic_vector (0 to 1 );
	f: out std_logic);
end WithSelect;

architecture Behavioral of WithSelect is
begin
	with a select
	f <= '1' when  "00",
		'1' when  "10",
		'1' when  "11",
		'0' when others;
end Behavioral;

