----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    08:29:11 11/24/2021 
-- Design Name: 
-- Module Name:    Lecccion3 - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity Lecccion3 is port(
	a,b: in std_logic;
	X: buffer std_logic_vector (1 downto 0);
	Z: buffer std_logic_vector (0 to 3));
end Lecccion3;

architecture Behavioral of Lecccion3 is
begin
	


end Behavioral;

